module ram_dp_4k (
    input           clk0_i,
    input           rst0_i,
    input   [ 13:0] addr0_i,
    input   [ 31:0] data0_i,
    input   [  3:0] wr0_i,
    input           clk1_i,
    input           rst1_i,
    input   [ 13:0] addr1_i,
    input   [ 31:0] data1_i,
    input   [  3:0] wr1_i,
    output  [ 31:0] data0_o,
    output  [ 31:0] data1_o
);

/* verilator lint_off MULTIDRIVEN */
reg [31:0]   ram [4095:0];
/* verilator lint_on MULTIDRIVEN */

initial $readmemh("../../../../ZYNQ_RISCV.sdk/app_test/app_test.txt", ram);

reg [31:0] ram_read0_q;
reg [31:0] ram_read1_q;

// Synchronous write
always @ (posedge clk0_i)
begin
    if (wr0_i[0])
        ram[addr0_i][7:0] <= data0_i[7:0];
    if (wr0_i[1])
        ram[addr0_i][15:8] <= data0_i[15:8];
    if (wr0_i[2])
        ram[addr0_i][23:16] <= data0_i[23:16];
    if (wr0_i[3])
        ram[addr0_i][31:24] <= data0_i[31:24];

    ram_read0_q <= ram[addr0_i];
end

always @ (posedge clk1_i)
begin
    if (wr1_i[0])
        ram[addr1_i][7:0] <= data1_i[7:0];
    if (wr1_i[1])
        ram[addr1_i][15:8] <= data1_i[15:8];
    if (wr1_i[2])
        ram[addr1_i][23:16] <= data1_i[23:16];
    if (wr1_i[3])
        ram[addr1_i][31:24] <= data1_i[31:24];

    ram_read1_q <= ram[addr1_i];
end

assign data0_o = ram_read0_q;
assign data1_o = ram_read1_q;


endmodule
